module greater (input [1:0] a, b,
                output      out);

   assign out = a > b;
endmodule
